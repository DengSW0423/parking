library ieee;
use ieee.std_logic_1164.all;

entity debouncer is
	port(
		clk_1000hz: in std_logic;
		btn_in: in std_logic;
		btn_out: out std_logic
	);
end debouncer;

architecture arch of debouncer is
begin
	process(clk_1000hz)
		variable count: integer range 0 to 25;
		variable btn_out_t: std_logic;
	begin
		if rising_edge(clk_1000hz) then
			if btn_in = '1' then
				if count = 25 then
					count := count;
				else
					count := count + 1;
				end if;
				
				if count = 24 then
					btn_out_t := '1';
				else
					btn_out_t := '0';
				end if;
			else
				count := 0;
			end if;
		end if; 
		
		btn_out <= btn_out_t;
	end process;
	
end arch;
