library ieee;
use ieee.std_logic_1164.all;
use work.my_package.all;

entity disp_driver is
	port(
		rst: in std_logic;
		clk_1000hz: in std_logic;
		clk_2hz: in std_logic;
		blinking: in boolean;
		numbers: in integer_array;
		disp: out std_logic_vector(6 downto 0);
		disp_switch: buffer bit_vector(5 downto 0)
	);
end disp_driver;

architecture arch of disp_driver is
	signal disp_left_0, disp_right_0: std_logic_vector(6 downto 0);
	signal disp_left_1, disp_right_1: std_logic_vector(6 downto 0);
	signal disp_left_2, disp_right_2: std_logic_vector(6 downto 0);
begin

	process(clk_1000hz, rst)
		variable disp_state: bit_vector(5 downto 0) := "111111";
	begin
		if rst = '1' then
			if disp_state = "111111" then
				disp_state := "011111";
			else
				disp_state := "111111";
			end if;
		elsif rising_edge(clk_1000hz) then
			if blinking and clk_2hz = '1' then
				disp_switch <= "111111";
			else
				disp_switch <= disp_state;
				case disp_state is
					when "011111" => disp <= disp_left_0;
					when "101111" => disp <= disp_right_0;
					when "110111" => disp <= disp_left_1;
					when "111011" => disp <= disp_right_1;
					when "111101" => disp <= disp_left_2;
					when "111110" => disp <= disp_right_2;
					when others => null;
				end case;
				disp_state := disp_state ror 1;
			end if;
		end if;
	end process;
	
	process(numbers(0))
	begin
		case numbers(0) is
			when 0 => disp_left_0 <= ZERO; disp_right_0 <= ZERO;
			when 1 => disp_left_0 <= ZERO; disp_right_0 <= ONE;
			when 2 => disp_left_0 <= ZERO; disp_right_0 <= TWO;
			when 3 => disp_left_0 <= ZERO; disp_right_0 <= THREE;
			when 4 => disp_left_0 <= ZERO; disp_right_0 <= FOUR;
			when 5 => disp_left_0 <= ZERO; disp_right_0 <= FIVE;
			when 6 => disp_left_0 <= ZERO; disp_right_0 <= SIX;
			when 7 => disp_left_0 <= ZERO; disp_right_0 <= SEVEN;
			when 8 => disp_left_0 <= ZERO; disp_right_0 <= EIGHT;
			when 9 => disp_left_0 <= ZERO; disp_right_0 <= NINE;
			when 10 => disp_left_0 <= ONE; disp_right_0 <= ZERO;
			when 11 => disp_left_0 <= ONE; disp_right_0 <= ONE;
			when 12 => disp_left_0 <= ONE; disp_right_0 <= TWO;
			when 13 => disp_left_0 <= ONE; disp_right_0 <= THREE;
			when 14 => disp_left_0 <= ONE; disp_right_0 <= FOUR;
			when 15 => disp_left_0 <= ONE; disp_right_0 <= FIVE;
			when 16 => disp_left_0 <= ONE; disp_right_0 <= SIX;
			when 17 => disp_left_0 <= ONE; disp_right_0 <= SEVEN;
			when 18 => disp_left_0 <= ONE; disp_right_0 <= EIGHT;
			when 19 => disp_left_0 <= ONE; disp_right_0 <= NINE;
			when 20 => disp_left_0 <= TWO; disp_right_0 <= ZERO;
			when 21 => disp_left_0 <= TWO; disp_right_0 <= ONE;
			when 22 => disp_left_0 <= TWO; disp_right_0 <= TWO;
			when 23 => disp_left_0 <= TWO; disp_right_0 <= THREE;
			when 24 => disp_left_0 <= TWO; disp_right_0 <= FOUR;
			when 25 => disp_left_0 <= TWO; disp_right_0 <= FIVE;
			when 26 => disp_left_0 <= TWO; disp_right_0 <= SIX;
			when 27 => disp_left_0 <= TWO; disp_right_0 <= SEVEN;
			when 28 => disp_left_0 <= TWO; disp_right_0 <= EIGHT;
			when 29 => disp_left_0 <= TWO; disp_right_0 <= NINE;
			when 30 => disp_left_0 <= THREE; disp_right_0 <= ZERO;
			when 31 => disp_left_0 <= THREE; disp_right_0 <= ONE;
			when 32 => disp_left_0 <= THREE; disp_right_0 <= TWO;
			when 33 => disp_left_0 <= THREE; disp_right_0 <= THREE;
			when 34 => disp_left_0 <= THREE; disp_right_0 <= FOUR;
			when 35 => disp_left_0 <= THREE; disp_right_0 <= FIVE;
			when 36 => disp_left_0 <= THREE; disp_right_0 <= SIX;
			when 37 => disp_left_0 <= THREE; disp_right_0 <= SEVEN;
			when 38 => disp_left_0 <= THREE; disp_right_0 <= EIGHT;
			when 39 => disp_left_0 <= THREE; disp_right_0 <= NINE;
			when 40 => disp_left_0 <= FOUR; disp_right_0 <= ZERO;
			when 41 => disp_left_0 <= FOUR; disp_right_0 <= ONE;
			when 42 => disp_left_0 <= FOUR; disp_right_0 <= TWO;
			when 43 => disp_left_0 <= FOUR; disp_right_0 <= THREE;
			when 44 => disp_left_0 <= FOUR; disp_right_0 <= FOUR;
			when 45 => disp_left_0 <= FOUR; disp_right_0 <= FIVE;
			when 46 => disp_left_0 <= FOUR; disp_right_0 <= SIX;
			when 47 => disp_left_0 <= FOUR; disp_right_0 <= SEVEN;
			when 48 => disp_left_0 <= FOUR; disp_right_0 <= EIGHT;
			when 49 => disp_left_0 <= FOUR; disp_right_0 <= NINE;
			when 50 => disp_left_0 <= FIVE; disp_right_0 <= ZERO;
			when 51 => disp_left_0 <= FIVE; disp_right_0 <= ONE;
			when 52 => disp_left_0 <= FIVE; disp_right_0 <= TWO;
			when 53 => disp_left_0 <= FIVE; disp_right_0 <= THREE;
			when 54 => disp_left_0 <= FIVE; disp_right_0 <= FOUR;
			when 55 => disp_left_0 <= FIVE; disp_right_0 <= FIVE;
			when 56 => disp_left_0 <= FIVE; disp_right_0 <= SIX;
			when 57 => disp_left_0 <= FIVE; disp_right_0 <= SEVEN;
			when 58 => disp_left_0 <= FIVE; disp_right_0 <= EIGHT;
			when 59 => disp_left_0 <= FIVE; disp_right_0 <= NINE;
			when 60 => disp_left_0 <= SIX; disp_right_0 <= ZERO;
			when 61 => disp_left_0 <= SIX; disp_right_0 <= ONE;
			when 62 => disp_left_0 <= SIX; disp_right_0 <= TWO;
			when 63 => disp_left_0 <= SIX; disp_right_0 <= THREE;
			when 64 => disp_left_0 <= SIX; disp_right_0 <= FOUR;
			when 65 => disp_left_0 <= SIX; disp_right_0 <= FIVE;
			when 66 => disp_left_0 <= SIX; disp_right_0 <= SIX;
			when 67 => disp_left_0 <= SIX; disp_right_0 <= SEVEN;
			when 68 => disp_left_0 <= SIX; disp_right_0 <= EIGHT;
			when 69 => disp_left_0 <= SIX; disp_right_0 <= NINE;
			when 70 => disp_left_0 <= SEVEN; disp_right_0 <= ZERO;
			when 71 => disp_left_0 <= SEVEN; disp_right_0 <= ONE;
			when 72 => disp_left_0 <= SEVEN; disp_right_0 <= TWO;
			when 73 => disp_left_0 <= SEVEN; disp_right_0 <= THREE;
			when 74 => disp_left_0 <= SEVEN; disp_right_0 <= FOUR;
			when 75 => disp_left_0 <= SEVEN; disp_right_0 <= FIVE;
			when 76 => disp_left_0 <= SEVEN; disp_right_0 <= SIX;
			when 77 => disp_left_0 <= SEVEN; disp_right_0 <= SEVEN;
			when 78 => disp_left_0 <= SEVEN; disp_right_0 <= EIGHT;
			when 79 => disp_left_0 <= SEVEN; disp_right_0 <= NINE;
			when 80 => disp_left_0 <= EIGHT; disp_right_0 <= ZERO;
			when 81 => disp_left_0 <= EIGHT; disp_right_0 <= ONE;
			when 82 => disp_left_0 <= EIGHT; disp_right_0 <= TWO;
			when 83 => disp_left_0 <= EIGHT; disp_right_0 <= THREE;
			when 84 => disp_left_0 <= EIGHT; disp_right_0 <= FOUR;
			when 85 => disp_left_0 <= EIGHT; disp_right_0 <= FIVE;
			when 86 => disp_left_0 <= EIGHT; disp_right_0 <= SIX;
			when 87 => disp_left_0 <= EIGHT; disp_right_0 <= SEVEN;
			when 88 => disp_left_0 <= EIGHT; disp_right_0 <= EIGHT;
			when 89 => disp_left_0 <= EIGHT; disp_right_0 <= NINE;
			when 90 => disp_left_0 <= NINE; disp_right_0 <= ZERO;
			when 91 => disp_left_0 <= NINE; disp_right_0 <= ONE;
			when 92 => disp_left_0 <= NINE; disp_right_0 <= TWO;
			when 93 => disp_left_0 <= NINE; disp_right_0 <= THREE;
			when 94 => disp_left_0 <= NINE; disp_right_0 <= FOUR;
			when 95 => disp_left_0 <= NINE; disp_right_0 <= FIVE;
			when 96 => disp_left_0 <= NINE; disp_right_0 <= SIX;
			when 97 => disp_left_0 <= NINE; disp_right_0 <= SEVEN;
			when 98 => disp_left_0 <= NINE; disp_right_0 <= EIGHT;
			when 99 => disp_left_0 <= NINE; disp_right_0 <= NINE;
			when others => null;
		end case;
	end process;
	
	process(numbers(1))
	begin
		case numbers(1) is
			when 0 => disp_left_1 <= ZERO; disp_right_1 <= ZERO;
			when 1 => disp_left_1 <= ZERO; disp_right_1 <= ONE;
			when 2 => disp_left_1 <= ZERO; disp_right_1 <= TWO;
			when 3 => disp_left_1 <= ZERO; disp_right_1 <= THREE;
			when 4 => disp_left_1 <= ZERO; disp_right_1 <= FOUR;
			when 5 => disp_left_1 <= ZERO; disp_right_1 <= FIVE;
			when 6 => disp_left_1 <= ZERO; disp_right_1 <= SIX;
			when 7 => disp_left_1 <= ZERO; disp_right_1 <= SEVEN;
			when 8 => disp_left_1 <= ZERO; disp_right_1 <= EIGHT;
			when 9 => disp_left_1 <= ZERO; disp_right_1 <= NINE;
			when 10 => disp_left_1 <= ONE; disp_right_1 <= ZERO;
			when 11 => disp_left_1 <= ONE; disp_right_1 <= ONE;
			when 12 => disp_left_1 <= ONE; disp_right_1 <= TWO;
			when 13 => disp_left_1 <= ONE; disp_right_1 <= THREE;
			when 14 => disp_left_1 <= ONE; disp_right_1 <= FOUR;
			when 15 => disp_left_1 <= ONE; disp_right_1 <= FIVE;
			when 16 => disp_left_1 <= ONE; disp_right_1 <= SIX;
			when 17 => disp_left_1 <= ONE; disp_right_1 <= SEVEN;
			when 18 => disp_left_1 <= ONE; disp_right_1 <= EIGHT;
			when 19 => disp_left_1 <= ONE; disp_right_1 <= NINE;
			when 20 => disp_left_1 <= TWO; disp_right_1 <= ZERO;
			when 21 => disp_left_1 <= TWO; disp_right_1 <= ONE;
			when 22 => disp_left_1 <= TWO; disp_right_1 <= TWO;
			when 23 => disp_left_1 <= TWO; disp_right_1 <= THREE;
			when 24 => disp_left_1 <= TWO; disp_right_1 <= FOUR;
			when 25 => disp_left_1 <= TWO; disp_right_1 <= FIVE;
			when 26 => disp_left_1 <= TWO; disp_right_1 <= SIX;
			when 27 => disp_left_1 <= TWO; disp_right_1 <= SEVEN;
			when 28 => disp_left_1 <= TWO; disp_right_1 <= EIGHT;
			when 29 => disp_left_1 <= TWO; disp_right_1 <= NINE;
			when 30 => disp_left_1 <= THREE; disp_right_1 <= ZERO;
			when 31 => disp_left_1 <= THREE; disp_right_1 <= ONE;
			when 32 => disp_left_1 <= THREE; disp_right_1 <= TWO;
			when 33 => disp_left_1 <= THREE; disp_right_1 <= THREE;
			when 34 => disp_left_1 <= THREE; disp_right_1 <= FOUR;
			when 35 => disp_left_1 <= THREE; disp_right_1 <= FIVE;
			when 36 => disp_left_1 <= THREE; disp_right_1 <= SIX;
			when 37 => disp_left_1 <= THREE; disp_right_1 <= SEVEN;
			when 38 => disp_left_1 <= THREE; disp_right_1 <= EIGHT;
			when 39 => disp_left_1 <= THREE; disp_right_1 <= NINE;
			when 40 => disp_left_1 <= FOUR; disp_right_1 <= ZERO;
			when 41 => disp_left_1 <= FOUR; disp_right_1 <= ONE;
			when 42 => disp_left_1 <= FOUR; disp_right_1 <= TWO;
			when 43 => disp_left_1 <= FOUR; disp_right_1 <= THREE;
			when 44 => disp_left_1 <= FOUR; disp_right_1 <= FOUR;
			when 45 => disp_left_1 <= FOUR; disp_right_1 <= FIVE;
			when 46 => disp_left_1 <= FOUR; disp_right_1 <= SIX;
			when 47 => disp_left_1 <= FOUR; disp_right_1 <= SEVEN;
			when 48 => disp_left_1 <= FOUR; disp_right_1 <= EIGHT;
			when 49 => disp_left_1 <= FOUR; disp_right_1 <= NINE;
			when 50 => disp_left_1 <= FIVE; disp_right_1 <= ZERO;
			when 51 => disp_left_1 <= FIVE; disp_right_1 <= ONE;
			when 52 => disp_left_1 <= FIVE; disp_right_1 <= TWO;
			when 53 => disp_left_1 <= FIVE; disp_right_1 <= THREE;
			when 54 => disp_left_1 <= FIVE; disp_right_1 <= FOUR;
			when 55 => disp_left_1 <= FIVE; disp_right_1 <= FIVE;
			when 56 => disp_left_1 <= FIVE; disp_right_1 <= SIX;
			when 57 => disp_left_1 <= FIVE; disp_right_1 <= SEVEN;
			when 58 => disp_left_1 <= FIVE; disp_right_1 <= EIGHT;
			when 59 => disp_left_1 <= FIVE; disp_right_1 <= NINE;
			when 60 => disp_left_1 <= SIX; disp_right_1 <= ZERO;
			when 61 => disp_left_1 <= SIX; disp_right_1 <= ONE;
			when 62 => disp_left_1 <= SIX; disp_right_1 <= TWO;
			when 63 => disp_left_1 <= SIX; disp_right_1 <= THREE;
			when 64 => disp_left_1 <= SIX; disp_right_1 <= FOUR;
			when 65 => disp_left_1 <= SIX; disp_right_1 <= FIVE;
			when 66 => disp_left_1 <= SIX; disp_right_1 <= SIX;
			when 67 => disp_left_1 <= SIX; disp_right_1 <= SEVEN;
			when 68 => disp_left_1 <= SIX; disp_right_1 <= EIGHT;
			when 69 => disp_left_1 <= SIX; disp_right_1 <= NINE;
			when 70 => disp_left_1 <= SEVEN; disp_right_1 <= ZERO;
			when 71 => disp_left_1 <= SEVEN; disp_right_1 <= ONE;
			when 72 => disp_left_1 <= SEVEN; disp_right_1 <= TWO;
			when 73 => disp_left_1 <= SEVEN; disp_right_1 <= THREE;
			when 74 => disp_left_1 <= SEVEN; disp_right_1 <= FOUR;
			when 75 => disp_left_1 <= SEVEN; disp_right_1 <= FIVE;
			when 76 => disp_left_1 <= SEVEN; disp_right_1 <= SIX;
			when 77 => disp_left_1 <= SEVEN; disp_right_1 <= SEVEN;
			when 78 => disp_left_1 <= SEVEN; disp_right_1 <= EIGHT;
			when 79 => disp_left_1 <= SEVEN; disp_right_1 <= NINE;
			when 80 => disp_left_1 <= EIGHT; disp_right_1 <= ZERO;
			when 81 => disp_left_1 <= EIGHT; disp_right_1 <= ONE;
			when 82 => disp_left_1 <= EIGHT; disp_right_1 <= TWO;
			when 83 => disp_left_1 <= EIGHT; disp_right_1 <= THREE;
			when 84 => disp_left_1 <= EIGHT; disp_right_1 <= FOUR;
			when 85 => disp_left_1 <= EIGHT; disp_right_1 <= FIVE;
			when 86 => disp_left_1 <= EIGHT; disp_right_1 <= SIX;
			when 87 => disp_left_1 <= EIGHT; disp_right_1 <= SEVEN;
			when 88 => disp_left_1 <= EIGHT; disp_right_1 <= EIGHT;
			when 89 => disp_left_1 <= EIGHT; disp_right_1 <= NINE;
			when 90 => disp_left_1 <= NINE; disp_right_1 <= ZERO;
			when 91 => disp_left_1 <= NINE; disp_right_1 <= ONE;
			when 92 => disp_left_1 <= NINE; disp_right_1 <= TWO;
			when 93 => disp_left_1 <= NINE; disp_right_1 <= THREE;
			when 94 => disp_left_1 <= NINE; disp_right_1 <= FOUR;
			when 95 => disp_left_1 <= NINE; disp_right_1 <= FIVE;
			when 96 => disp_left_1 <= NINE; disp_right_1 <= SIX;
			when 97 => disp_left_1 <= NINE; disp_right_1 <= SEVEN;
			when 98 => disp_left_1 <= NINE; disp_right_1 <= EIGHT;
			when 99 => disp_left_1 <= NINE; disp_right_1 <= NINE;
			when others => null;
		end case;
	end process;
	
	process(numbers(2))
	begin
		case numbers(2) is
			when 0 => disp_left_2 <= ZERO; disp_right_2 <= ZERO;
			when 1 => disp_left_2 <= ZERO; disp_right_2 <= ONE;
			when 2 => disp_left_2 <= ZERO; disp_right_2 <= TWO;
			when 3 => disp_left_2 <= ZERO; disp_right_2 <= THREE;
			when 4 => disp_left_2 <= ZERO; disp_right_2 <= FOUR;
			when 5 => disp_left_2 <= ZERO; disp_right_2 <= FIVE;
			when 6 => disp_left_2 <= ZERO; disp_right_2 <= SIX;
			when 7 => disp_left_2 <= ZERO; disp_right_2 <= SEVEN;
			when 8 => disp_left_2 <= ZERO; disp_right_2 <= EIGHT;
			when 9 => disp_left_2 <= ZERO; disp_right_2 <= NINE;
			when 10 => disp_left_2 <= ONE; disp_right_2 <= ZERO;
			when 11 => disp_left_2 <= ONE; disp_right_2 <= ONE;
			when 12 => disp_left_2 <= ONE; disp_right_2 <= TWO;
			when 13 => disp_left_2 <= ONE; disp_right_2 <= THREE;
			when 14 => disp_left_2 <= ONE; disp_right_2 <= FOUR;
			when 15 => disp_left_2 <= ONE; disp_right_2 <= FIVE;
			when 16 => disp_left_2 <= ONE; disp_right_2 <= SIX;
			when 17 => disp_left_2 <= ONE; disp_right_2 <= SEVEN;
			when 18 => disp_left_2 <= ONE; disp_right_2 <= EIGHT;
			when 19 => disp_left_2 <= ONE; disp_right_2 <= NINE;
			when 20 => disp_left_2 <= TWO; disp_right_2 <= ZERO;
			when 21 => disp_left_2 <= TWO; disp_right_2 <= ONE;
			when 22 => disp_left_2 <= TWO; disp_right_2 <= TWO;
			when 23 => disp_left_2 <= TWO; disp_right_2 <= THREE;
			when 24 => disp_left_2 <= TWO; disp_right_2 <= FOUR;
			when 25 => disp_left_2 <= TWO; disp_right_2 <= FIVE;
			when 26 => disp_left_2 <= TWO; disp_right_2 <= SIX;
			when 27 => disp_left_2 <= TWO; disp_right_2 <= SEVEN;
			when 28 => disp_left_2 <= TWO; disp_right_2 <= EIGHT;
			when 29 => disp_left_2 <= TWO; disp_right_2 <= NINE;
			when 30 => disp_left_2 <= THREE; disp_right_2 <= ZERO;
			when 31 => disp_left_2 <= THREE; disp_right_2 <= ONE;
			when 32 => disp_left_2 <= THREE; disp_right_2 <= TWO;
			when 33 => disp_left_2 <= THREE; disp_right_2 <= THREE;
			when 34 => disp_left_2 <= THREE; disp_right_2 <= FOUR;
			when 35 => disp_left_2 <= THREE; disp_right_2 <= FIVE;
			when 36 => disp_left_2 <= THREE; disp_right_2 <= SIX;
			when 37 => disp_left_2 <= THREE; disp_right_2 <= SEVEN;
			when 38 => disp_left_2 <= THREE; disp_right_2 <= EIGHT;
			when 39 => disp_left_2 <= THREE; disp_right_2 <= NINE;
			when 40 => disp_left_2 <= FOUR; disp_right_2 <= ZERO;
			when 41 => disp_left_2 <= FOUR; disp_right_2 <= ONE;
			when 42 => disp_left_2 <= FOUR; disp_right_2 <= TWO;
			when 43 => disp_left_2 <= FOUR; disp_right_2 <= THREE;
			when 44 => disp_left_2 <= FOUR; disp_right_2 <= FOUR;
			when 45 => disp_left_2 <= FOUR; disp_right_2 <= FIVE;
			when 46 => disp_left_2 <= FOUR; disp_right_2 <= SIX;
			when 47 => disp_left_2 <= FOUR; disp_right_2 <= SEVEN;
			when 48 => disp_left_2 <= FOUR; disp_right_2 <= EIGHT;
			when 49 => disp_left_2 <= FOUR; disp_right_2 <= NINE;
			when 50 => disp_left_2 <= FIVE; disp_right_2 <= ZERO;
			when 51 => disp_left_2 <= FIVE; disp_right_2 <= ONE;
			when 52 => disp_left_2 <= FIVE; disp_right_2 <= TWO;
			when 53 => disp_left_2 <= FIVE; disp_right_2 <= THREE;
			when 54 => disp_left_2 <= FIVE; disp_right_2 <= FOUR;
			when 55 => disp_left_2 <= FIVE; disp_right_2 <= FIVE;
			when 56 => disp_left_2 <= FIVE; disp_right_2 <= SIX;
			when 57 => disp_left_2 <= FIVE; disp_right_2 <= SEVEN;
			when 58 => disp_left_2 <= FIVE; disp_right_2 <= EIGHT;
			when 59 => disp_left_2 <= FIVE; disp_right_2 <= NINE;
			when 60 => disp_left_2 <= SIX; disp_right_2 <= ZERO;
			when 61 => disp_left_2 <= SIX; disp_right_2 <= ONE;
			when 62 => disp_left_2 <= SIX; disp_right_2 <= TWO;
			when 63 => disp_left_2 <= SIX; disp_right_2 <= THREE;
			when 64 => disp_left_2 <= SIX; disp_right_2 <= FOUR;
			when 65 => disp_left_2 <= SIX; disp_right_2 <= FIVE;
			when 66 => disp_left_2 <= SIX; disp_right_2 <= SIX;
			when 67 => disp_left_2 <= SIX; disp_right_2 <= SEVEN;
			when 68 => disp_left_2 <= SIX; disp_right_2 <= EIGHT;
			when 69 => disp_left_2 <= SIX; disp_right_2 <= NINE;
			when 70 => disp_left_2 <= SEVEN; disp_right_2 <= ZERO;
			when 71 => disp_left_2 <= SEVEN; disp_right_2 <= ONE;
			when 72 => disp_left_2 <= SEVEN; disp_right_2 <= TWO;
			when 73 => disp_left_2 <= SEVEN; disp_right_2 <= THREE;
			when 74 => disp_left_2 <= SEVEN; disp_right_2 <= FOUR;
			when 75 => disp_left_2 <= SEVEN; disp_right_2 <= FIVE;
			when 76 => disp_left_2 <= SEVEN; disp_right_2 <= SIX;
			when 77 => disp_left_2 <= SEVEN; disp_right_2 <= SEVEN;
			when 78 => disp_left_2 <= SEVEN; disp_right_2 <= EIGHT;
			when 79 => disp_left_2 <= SEVEN; disp_right_2 <= NINE;
			when 80 => disp_left_2 <= EIGHT; disp_right_2 <= ZERO;
			when 81 => disp_left_2 <= EIGHT; disp_right_2 <= ONE;
			when 82 => disp_left_2 <= EIGHT; disp_right_2 <= TWO;
			when 83 => disp_left_2 <= EIGHT; disp_right_2 <= THREE;
			when 84 => disp_left_2 <= EIGHT; disp_right_2 <= FOUR;
			when 85 => disp_left_2 <= EIGHT; disp_right_2 <= FIVE;
			when 86 => disp_left_2 <= EIGHT; disp_right_2 <= SIX;
			when 87 => disp_left_2 <= EIGHT; disp_right_2 <= SEVEN;
			when 88 => disp_left_2 <= EIGHT; disp_right_2 <= EIGHT;
			when 89 => disp_left_2 <= EIGHT; disp_right_2 <= NINE;
			when 90 => disp_left_2 <= NINE; disp_right_2 <= ZERO;
			when 91 => disp_left_2 <= NINE; disp_right_2 <= ONE;
			when 92 => disp_left_2 <= NINE; disp_right_2 <= TWO;
			when 93 => disp_left_2 <= NINE; disp_right_2 <= THREE;
			when 94 => disp_left_2 <= NINE; disp_right_2 <= FOUR;
			when 95 => disp_left_2 <= NINE; disp_right_2 <= FIVE;
			when 96 => disp_left_2 <= NINE; disp_right_2 <= SIX;
			when 97 => disp_left_2 <= NINE; disp_right_2 <= SEVEN;
			when 98 => disp_left_2 <= NINE; disp_right_2 <= EIGHT;
			when 99 => disp_left_2 <= NINE; disp_right_2 <= NINE;
			when others => null;
		end case;
	end process;
end arch;
