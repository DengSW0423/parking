library ieee;
use ieee.std_logic_1164.all;

entity initializer is
	port(
	
	);
end initializer;

architecture arch of initializer is

begin

end arch;
